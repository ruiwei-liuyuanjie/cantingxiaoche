////////////////////////////////////////////////////////////////////////////////
// SubModule main
// Created   2017/4/24 21:43:17
////////////////////////////////////////////////////////////////////////////////

module main (PCIE_CTX, PCIE_CRX, SONAR_TRIG4, MOTO_L_PWM, MOTO_R_PWM, SONAR_TRIG3, SONAR_TRIG2, SONAR_TRIG1, SONAR_ECHO4, SONAR_ECHO3, SONAR_ECHO2, SONAR_ECHO1, BATT_FAULT, BATT_CHRG, BATT_READY, HOME_IR_R3, HOME_IR_R2, HOME_IR_R1, GROUND_DETECT_R, MOTO_LB_EN, MOTO_RB_EN, MOTO_RF_EN, MOTO_LI_MONITOR, MOTO_LF_EN, ENCODER_SENSOR_L, ENCODER_SENSOR_R, GROUND_DETECT_L, PC10_RX, PC10_TX, PCIE_nCCMD, MOTTOM_IR_E, MOTO_RI_MONITOR, BOTTOM_IR_R3, BATT_MONITOR, BOTTOM_IR_R1, BOTTOM_IR_R2, CURRENT_SET, BUMP_DETECT_R, DCCHARGE_DETECT, HOCHARGE_DETECT, BUMP_DETECT_L, PCIE_CBUSY, BATT_DETECT, BOTTOM_IR_R4, UART2_RX_PA3, UART2_TX_PA2, CHARGE_PWM);

output PCIE_CTX;
output PCIE_CRX;
output SONAR_TRIG4;
output MOTO_L_PWM;
output MOTO_R_PWM;
output SONAR_TRIG3;
output SONAR_TRIG2;
output SONAR_TRIG1;
output SONAR_ECHO4;
output SONAR_ECHO3;
output SONAR_ECHO2;
output SONAR_ECHO1;
output BATT_FAULT;
output BATT_CHRG;
output BATT_READY;
output HOME_IR_R3;
output HOME_IR_R2;
output HOME_IR_R1;
output GROUND_DETECT_R;
output MOTO_LB_EN;
output MOTO_RB_EN;
output MOTO_RF_EN;
output MOTO_LI_MONITOR;
output MOTO_LF_EN;
output ENCODER_SENSOR_L;
output ENCODER_SENSOR_R;
output GROUND_DETECT_L;
output PC10_RX;
output PC10_TX;
output PCIE_nCCMD;
output MOTTOM_IR_E;
output MOTO_RI_MONITOR;
output BOTTOM_IR_R3;
output BATT_MONITOR;
output BOTTOM_IR_R1;
output BOTTOM_IR_R2;
output CURRENT_SET;
output BUMP_DETECT_R;
output DCCHARGE_DETECT;
output HOCHARGE_DETECT;
output BUMP_DETECT_L;
output PCIE_CBUSY;
output BATT_DETECT;
output BOTTOM_IR_R4;
output UART2_RX_PA3;
output UART2_TX_PA2;
output CHARGE_PWM;


endmodule
////////////////////////////////////////////////////////////////////////////////
